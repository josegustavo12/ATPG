`timescale 1ns/1ps
module tb;

  reg N1;
  reg N18;
  reg N35;
  reg N52;
  reg N69;
  reg N86;
  reg N103;
  reg N120;
  reg N137;
  reg N154;
  reg N171;
  reg N188;
  reg N205;
  reg N222;
  reg N239;
  reg N256;
  reg N273;
  reg N290;
  reg N307;
  reg N324;
  reg N341;
  reg N358;
  reg N375;
  reg N392;
  reg N409;
  reg N426;
  reg N443;
  reg N460;
  reg N477;
  reg N494;
  reg N511;
  reg N528;
  wire N545;
  wire N1581;
  wire N1901;
  wire N2223;
  wire N2548;
  wire N2877;
  wire N3211;
  wire N3552;
  wire N3895;
  wire N4241;
  wire N4591;
  wire N4946;
  wire N5308;
  wire N5672;
  wire N5971;
  wire N6123;
  wire N6150;
  wire N6160;
  wire N6170;
  wire N6180;
  wire N6190;
  wire N6200;
  wire N6210;
  wire N6220;
  wire N6230;
  wire N6240;
  wire N6250;
  wire N6260;
  wire N6270;
  wire N6280;
  wire N6287;
  wire N6288;

  c6288 uut (.N1(N1), .N18(N18), .N35(N35), .N52(N52), .N69(N69), .N86(N86), .N103(N103), .N120(N120), .N137(N137), .N154(N154), .N171(N171), .N188(N188), .N205(N205), .N222(N222), .N239(N239), .N256(N256), .N273(N273), .N290(N290), .N307(N307), .N324(N324), .N341(N341), .N358(N358), .N375(N375), .N392(N392), .N409(N409), .N426(N426), .N443(N443), .N460(N460), .N477(N477), .N494(N494), .N511(N511), .N528(N528), .N545(N545), .N1581(N1581), .N1901(N1901), .N2223(N2223), .N2548(N2548), .N2877(N2877), .N3211(N3211), .N3552(N3552), .N3895(N3895), .N4241(N4241), .N4591(N4591), .N4946(N4946), .N5308(N5308), .N5672(N5672), .N5971(N5971), .N6123(N6123), .N6150(N6150), .N6160(N6160), .N6170(N6170), .N6180(N6180), .N6190(N6190), .N6200(N6200), .N6210(N6210), .N6220(N6220), .N6230(N6230), .N6240(N6240), .N6250(N6250), .N6260(N6260), .N6270(N6270), .N6280(N6280), .N6287(N6287), .N6288(N6288));
  initial begin
    // Aplicando vetor 1
    N1 = 0;
    N18 = 0;
    N35 = 0;
    N52 = 1;
    N69 = 0;
    N86 = 0;
    N103 = 0;
    N120 = 0;
    N137 = 1;
    N154 = 0;
    N171 = 0;
    N188 = 0;
    N205 = 0;
    N222 = 1;
    N239 = 1;
    N256 = 0;
    N273 = 0;
    N290 = 0;
    N307 = 1;
    N324 = 1;
    N341 = 1;
    N358 = 0;
    N375 = 1;
    N392 = 1;
    N409 = 0;
    N426 = 0;
    N443 = 0;
    N460 = 0;
    N477 = 0;
    N494 = 0;
    N511 = 1;
    N528 = 0;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("1. OUTPUT: N545 = %b", N545);
    $display("1. OUTPUT: N1581 = %b", N1581);
    $display("1. OUTPUT: N1901 = %b", N1901);
    $display("1. OUTPUT: N2223 = %b", N2223);
    $display("1. OUTPUT: N2548 = %b", N2548);
    $display("1. OUTPUT: N2877 = %b", N2877);
    $display("1. OUTPUT: N3211 = %b", N3211);
    $display("1. OUTPUT: N3552 = %b", N3552);
    $display("1. OUTPUT: N3895 = %b", N3895);
    $display("1. OUTPUT: N4241 = %b", N4241);
    $display("1. OUTPUT: N4591 = %b", N4591);
    $display("1. OUTPUT: N4946 = %b", N4946);
    $display("1. OUTPUT: N5308 = %b", N5308);
    $display("1. OUTPUT: N5672 = %b", N5672);
    $display("1. OUTPUT: N5971 = %b", N5971);
    $display("1. OUTPUT: N6123 = %b", N6123);
    $display("1. OUTPUT: N6150 = %b", N6150);
    $display("1. OUTPUT: N6160 = %b", N6160);
    $display("1. OUTPUT: N6170 = %b", N6170);
    $display("1. OUTPUT: N6180 = %b", N6180);
    $display("1. OUTPUT: N6190 = %b", N6190);
    $display("1. OUTPUT: N6200 = %b", N6200);
    $display("1. OUTPUT: N6210 = %b", N6210);
    $display("1. OUTPUT: N6220 = %b", N6220);
    $display("1. OUTPUT: N6230 = %b", N6230);
    $display("1. OUTPUT: N6240 = %b", N6240);
    $display("1. OUTPUT: N6250 = %b", N6250);
    $display("1. OUTPUT: N6260 = %b", N6260);
    $display("1. OUTPUT: N6270 = %b", N6270);
    $display("1. OUTPUT: N6280 = %b", N6280);
    $display("1. OUTPUT: N6287 = %b", N6287);
    $display("1. OUTPUT: N6288 = %b", N6288);

    // Aplicando vetor 2
    N1 = 0;
    N18 = 0;
    N35 = 1;
    N52 = 1;
    N69 = 0;
    N86 = 0;
    N103 = 0;
    N120 = 1;
    N137 = 0;
    N154 = 1;
    N171 = 1;
    N188 = 0;
    N205 = 0;
    N222 = 0;
    N239 = 1;
    N256 = 1;
    N273 = 0;
    N290 = 1;
    N307 = 0;
    N324 = 1;
    N341 = 1;
    N358 = 1;
    N375 = 1;
    N392 = 1;
    N409 = 1;
    N426 = 1;
    N443 = 1;
    N460 = 0;
    N477 = 1;
    N494 = 1;
    N511 = 0;
    N528 = 0;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("2. OUTPUT: N545 = %b", N545);
    $display("2. OUTPUT: N1581 = %b", N1581);
    $display("2. OUTPUT: N1901 = %b", N1901);
    $display("2. OUTPUT: N2223 = %b", N2223);
    $display("2. OUTPUT: N2548 = %b", N2548);
    $display("2. OUTPUT: N2877 = %b", N2877);
    $display("2. OUTPUT: N3211 = %b", N3211);
    $display("2. OUTPUT: N3552 = %b", N3552);
    $display("2. OUTPUT: N3895 = %b", N3895);
    $display("2. OUTPUT: N4241 = %b", N4241);
    $display("2. OUTPUT: N4591 = %b", N4591);
    $display("2. OUTPUT: N4946 = %b", N4946);
    $display("2. OUTPUT: N5308 = %b", N5308);
    $display("2. OUTPUT: N5672 = %b", N5672);
    $display("2. OUTPUT: N5971 = %b", N5971);
    $display("2. OUTPUT: N6123 = %b", N6123);
    $display("2. OUTPUT: N6150 = %b", N6150);
    $display("2. OUTPUT: N6160 = %b", N6160);
    $display("2. OUTPUT: N6170 = %b", N6170);
    $display("2. OUTPUT: N6180 = %b", N6180);
    $display("2. OUTPUT: N6190 = %b", N6190);
    $display("2. OUTPUT: N6200 = %b", N6200);
    $display("2. OUTPUT: N6210 = %b", N6210);
    $display("2. OUTPUT: N6220 = %b", N6220);
    $display("2. OUTPUT: N6230 = %b", N6230);
    $display("2. OUTPUT: N6240 = %b", N6240);
    $display("2. OUTPUT: N6250 = %b", N6250);
    $display("2. OUTPUT: N6260 = %b", N6260);
    $display("2. OUTPUT: N6270 = %b", N6270);
    $display("2. OUTPUT: N6280 = %b", N6280);
    $display("2. OUTPUT: N6287 = %b", N6287);
    $display("2. OUTPUT: N6288 = %b", N6288);

    // Aplicando vetor 3
    N1 = 1;
    N18 = 1;
    N35 = 0;
    N52 = 0;
    N69 = 0;
    N86 = 1;
    N103 = 1;
    N120 = 0;
    N137 = 0;
    N154 = 1;
    N171 = 1;
    N188 = 1;
    N205 = 0;
    N222 = 1;
    N239 = 1;
    N256 = 1;
    N273 = 0;
    N290 = 1;
    N307 = 1;
    N324 = 1;
    N341 = 0;
    N358 = 1;
    N375 = 0;
    N392 = 1;
    N409 = 1;
    N426 = 0;
    N443 = 0;
    N460 = 1;
    N477 = 0;
    N494 = 1;
    N511 = 1;
    N528 = 1;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("3. OUTPUT: N545 = %b", N545);
    $display("3. OUTPUT: N1581 = %b", N1581);
    $display("3. OUTPUT: N1901 = %b", N1901);
    $display("3. OUTPUT: N2223 = %b", N2223);
    $display("3. OUTPUT: N2548 = %b", N2548);
    $display("3. OUTPUT: N2877 = %b", N2877);
    $display("3. OUTPUT: N3211 = %b", N3211);
    $display("3. OUTPUT: N3552 = %b", N3552);
    $display("3. OUTPUT: N3895 = %b", N3895);
    $display("3. OUTPUT: N4241 = %b", N4241);
    $display("3. OUTPUT: N4591 = %b", N4591);
    $display("3. OUTPUT: N4946 = %b", N4946);
    $display("3. OUTPUT: N5308 = %b", N5308);
    $display("3. OUTPUT: N5672 = %b", N5672);
    $display("3. OUTPUT: N5971 = %b", N5971);
    $display("3. OUTPUT: N6123 = %b", N6123);
    $display("3. OUTPUT: N6150 = %b", N6150);
    $display("3. OUTPUT: N6160 = %b", N6160);
    $display("3. OUTPUT: N6170 = %b", N6170);
    $display("3. OUTPUT: N6180 = %b", N6180);
    $display("3. OUTPUT: N6190 = %b", N6190);
    $display("3. OUTPUT: N6200 = %b", N6200);
    $display("3. OUTPUT: N6210 = %b", N6210);
    $display("3. OUTPUT: N6220 = %b", N6220);
    $display("3. OUTPUT: N6230 = %b", N6230);
    $display("3. OUTPUT: N6240 = %b", N6240);
    $display("3. OUTPUT: N6250 = %b", N6250);
    $display("3. OUTPUT: N6260 = %b", N6260);
    $display("3. OUTPUT: N6270 = %b", N6270);
    $display("3. OUTPUT: N6280 = %b", N6280);
    $display("3. OUTPUT: N6287 = %b", N6287);
    $display("3. OUTPUT: N6288 = %b", N6288);

    // Aplicando vetor 4
    N1 = 0;
    N18 = 0;
    N35 = 1;
    N52 = 1;
    N69 = 1;
    N86 = 0;
    N103 = 1;
    N120 = 1;
    N137 = 1;
    N154 = 0;
    N171 = 0;
    N188 = 0;
    N205 = 0;
    N222 = 0;
    N239 = 0;
    N256 = 0;
    N273 = 0;
    N290 = 1;
    N307 = 0;
    N324 = 1;
    N341 = 1;
    N358 = 1;
    N375 = 0;
    N392 = 1;
    N409 = 0;
    N426 = 1;
    N443 = 1;
    N460 = 0;
    N477 = 1;
    N494 = 0;
    N511 = 0;
    N528 = 1;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("4. OUTPUT: N545 = %b", N545);
    $display("4. OUTPUT: N1581 = %b", N1581);
    $display("4. OUTPUT: N1901 = %b", N1901);
    $display("4. OUTPUT: N2223 = %b", N2223);
    $display("4. OUTPUT: N2548 = %b", N2548);
    $display("4. OUTPUT: N2877 = %b", N2877);
    $display("4. OUTPUT: N3211 = %b", N3211);
    $display("4. OUTPUT: N3552 = %b", N3552);
    $display("4. OUTPUT: N3895 = %b", N3895);
    $display("4. OUTPUT: N4241 = %b", N4241);
    $display("4. OUTPUT: N4591 = %b", N4591);
    $display("4. OUTPUT: N4946 = %b", N4946);
    $display("4. OUTPUT: N5308 = %b", N5308);
    $display("4. OUTPUT: N5672 = %b", N5672);
    $display("4. OUTPUT: N5971 = %b", N5971);
    $display("4. OUTPUT: N6123 = %b", N6123);
    $display("4. OUTPUT: N6150 = %b", N6150);
    $display("4. OUTPUT: N6160 = %b", N6160);
    $display("4. OUTPUT: N6170 = %b", N6170);
    $display("4. OUTPUT: N6180 = %b", N6180);
    $display("4. OUTPUT: N6190 = %b", N6190);
    $display("4. OUTPUT: N6200 = %b", N6200);
    $display("4. OUTPUT: N6210 = %b", N6210);
    $display("4. OUTPUT: N6220 = %b", N6220);
    $display("4. OUTPUT: N6230 = %b", N6230);
    $display("4. OUTPUT: N6240 = %b", N6240);
    $display("4. OUTPUT: N6250 = %b", N6250);
    $display("4. OUTPUT: N6260 = %b", N6260);
    $display("4. OUTPUT: N6270 = %b", N6270);
    $display("4. OUTPUT: N6280 = %b", N6280);
    $display("4. OUTPUT: N6287 = %b", N6287);
    $display("4. OUTPUT: N6288 = %b", N6288);

    // Aplicando vetor 5
    N1 = 1;
    N18 = 1;
    N35 = 1;
    N52 = 0;
    N69 = 0;
    N86 = 0;
    N103 = 1;
    N120 = 1;
    N137 = 1;
    N154 = 0;
    N171 = 0;
    N188 = 0;
    N205 = 0;
    N222 = 1;
    N239 = 0;
    N256 = 0;
    N273 = 1;
    N290 = 1;
    N307 = 0;
    N324 = 1;
    N341 = 1;
    N358 = 1;
    N375 = 1;
    N392 = 1;
    N409 = 1;
    N426 = 1;
    N443 = 1;
    N460 = 1;
    N477 = 0;
    N494 = 1;
    N511 = 1;
    N528 = 1;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("5. OUTPUT: N545 = %b", N545);
    $display("5. OUTPUT: N1581 = %b", N1581);
    $display("5. OUTPUT: N1901 = %b", N1901);
    $display("5. OUTPUT: N2223 = %b", N2223);
    $display("5. OUTPUT: N2548 = %b", N2548);
    $display("5. OUTPUT: N2877 = %b", N2877);
    $display("5. OUTPUT: N3211 = %b", N3211);
    $display("5. OUTPUT: N3552 = %b", N3552);
    $display("5. OUTPUT: N3895 = %b", N3895);
    $display("5. OUTPUT: N4241 = %b", N4241);
    $display("5. OUTPUT: N4591 = %b", N4591);
    $display("5. OUTPUT: N4946 = %b", N4946);
    $display("5. OUTPUT: N5308 = %b", N5308);
    $display("5. OUTPUT: N5672 = %b", N5672);
    $display("5. OUTPUT: N5971 = %b", N5971);
    $display("5. OUTPUT: N6123 = %b", N6123);
    $display("5. OUTPUT: N6150 = %b", N6150);
    $display("5. OUTPUT: N6160 = %b", N6160);
    $display("5. OUTPUT: N6170 = %b", N6170);
    $display("5. OUTPUT: N6180 = %b", N6180);
    $display("5. OUTPUT: N6190 = %b", N6190);
    $display("5. OUTPUT: N6200 = %b", N6200);
    $display("5. OUTPUT: N6210 = %b", N6210);
    $display("5. OUTPUT: N6220 = %b", N6220);
    $display("5. OUTPUT: N6230 = %b", N6230);
    $display("5. OUTPUT: N6240 = %b", N6240);
    $display("5. OUTPUT: N6250 = %b", N6250);
    $display("5. OUTPUT: N6260 = %b", N6260);
    $display("5. OUTPUT: N6270 = %b", N6270);
    $display("5. OUTPUT: N6280 = %b", N6280);
    $display("5. OUTPUT: N6287 = %b", N6287);
    $display("5. OUTPUT: N6288 = %b", N6288);

    // Aplicando vetor 6
    N1 = 0;
    N18 = 1;
    N35 = 0;
    N52 = 1;
    N69 = 0;
    N86 = 0;
    N103 = 0;
    N120 = 1;
    N137 = 0;
    N154 = 1;
    N171 = 1;
    N188 = 0;
    N205 = 0;
    N222 = 1;
    N239 = 0;
    N256 = 1;
    N273 = 1;
    N290 = 1;
    N307 = 0;
    N324 = 0;
    N341 = 0;
    N358 = 0;
    N375 = 0;
    N392 = 0;
    N409 = 1;
    N426 = 1;
    N443 = 1;
    N460 = 1;
    N477 = 1;
    N494 = 1;
    N511 = 1;
    N528 = 1;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("6. OUTPUT: N545 = %b", N545);
    $display("6. OUTPUT: N1581 = %b", N1581);
    $display("6. OUTPUT: N1901 = %b", N1901);
    $display("6. OUTPUT: N2223 = %b", N2223);
    $display("6. OUTPUT: N2548 = %b", N2548);
    $display("6. OUTPUT: N2877 = %b", N2877);
    $display("6. OUTPUT: N3211 = %b", N3211);
    $display("6. OUTPUT: N3552 = %b", N3552);
    $display("6. OUTPUT: N3895 = %b", N3895);
    $display("6. OUTPUT: N4241 = %b", N4241);
    $display("6. OUTPUT: N4591 = %b", N4591);
    $display("6. OUTPUT: N4946 = %b", N4946);
    $display("6. OUTPUT: N5308 = %b", N5308);
    $display("6. OUTPUT: N5672 = %b", N5672);
    $display("6. OUTPUT: N5971 = %b", N5971);
    $display("6. OUTPUT: N6123 = %b", N6123);
    $display("6. OUTPUT: N6150 = %b", N6150);
    $display("6. OUTPUT: N6160 = %b", N6160);
    $display("6. OUTPUT: N6170 = %b", N6170);
    $display("6. OUTPUT: N6180 = %b", N6180);
    $display("6. OUTPUT: N6190 = %b", N6190);
    $display("6. OUTPUT: N6200 = %b", N6200);
    $display("6. OUTPUT: N6210 = %b", N6210);
    $display("6. OUTPUT: N6220 = %b", N6220);
    $display("6. OUTPUT: N6230 = %b", N6230);
    $display("6. OUTPUT: N6240 = %b", N6240);
    $display("6. OUTPUT: N6250 = %b", N6250);
    $display("6. OUTPUT: N6260 = %b", N6260);
    $display("6. OUTPUT: N6270 = %b", N6270);
    $display("6. OUTPUT: N6280 = %b", N6280);
    $display("6. OUTPUT: N6287 = %b", N6287);
    $display("6. OUTPUT: N6288 = %b", N6288);

    // Aplicando vetor 7
    N1 = 1;
    N18 = 0;
    N35 = 0;
    N52 = 0;
    N69 = 1;
    N86 = 1;
    N103 = 0;
    N120 = 1;
    N137 = 0;
    N154 = 0;
    N171 = 0;
    N188 = 0;
    N205 = 0;
    N222 = 0;
    N239 = 0;
    N256 = 1;
    N273 = 1;
    N290 = 0;
    N307 = 0;
    N324 = 1;
    N341 = 1;
    N358 = 1;
    N375 = 0;
    N392 = 0;
    N409 = 1;
    N426 = 1;
    N443 = 0;
    N460 = 1;
    N477 = 1;
    N494 = 1;
    N511 = 0;
    N528 = 0;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("7. OUTPUT: N545 = %b", N545);
    $display("7. OUTPUT: N1581 = %b", N1581);
    $display("7. OUTPUT: N1901 = %b", N1901);
    $display("7. OUTPUT: N2223 = %b", N2223);
    $display("7. OUTPUT: N2548 = %b", N2548);
    $display("7. OUTPUT: N2877 = %b", N2877);
    $display("7. OUTPUT: N3211 = %b", N3211);
    $display("7. OUTPUT: N3552 = %b", N3552);
    $display("7. OUTPUT: N3895 = %b", N3895);
    $display("7. OUTPUT: N4241 = %b", N4241);
    $display("7. OUTPUT: N4591 = %b", N4591);
    $display("7. OUTPUT: N4946 = %b", N4946);
    $display("7. OUTPUT: N5308 = %b", N5308);
    $display("7. OUTPUT: N5672 = %b", N5672);
    $display("7. OUTPUT: N5971 = %b", N5971);
    $display("7. OUTPUT: N6123 = %b", N6123);
    $display("7. OUTPUT: N6150 = %b", N6150);
    $display("7. OUTPUT: N6160 = %b", N6160);
    $display("7. OUTPUT: N6170 = %b", N6170);
    $display("7. OUTPUT: N6180 = %b", N6180);
    $display("7. OUTPUT: N6190 = %b", N6190);
    $display("7. OUTPUT: N6200 = %b", N6200);
    $display("7. OUTPUT: N6210 = %b", N6210);
    $display("7. OUTPUT: N6220 = %b", N6220);
    $display("7. OUTPUT: N6230 = %b", N6230);
    $display("7. OUTPUT: N6240 = %b", N6240);
    $display("7. OUTPUT: N6250 = %b", N6250);
    $display("7. OUTPUT: N6260 = %b", N6260);
    $display("7. OUTPUT: N6270 = %b", N6270);
    $display("7. OUTPUT: N6280 = %b", N6280);
    $display("7. OUTPUT: N6287 = %b", N6287);
    $display("7. OUTPUT: N6288 = %b", N6288);

    // Aplicando vetor 8
    N1 = 1;
    N18 = 0;
    N35 = 1;
    N52 = 1;
    N69 = 1;
    N86 = 0;
    N103 = 1;
    N120 = 1;
    N137 = 1;
    N154 = 1;
    N171 = 1;
    N188 = 1;
    N205 = 0;
    N222 = 1;
    N239 = 0;
    N256 = 1;
    N273 = 0;
    N290 = 1;
    N307 = 1;
    N324 = 0;
    N341 = 1;
    N358 = 1;
    N375 = 1;
    N392 = 0;
    N409 = 0;
    N426 = 1;
    N443 = 1;
    N460 = 1;
    N477 = 0;
    N494 = 1;
    N511 = 0;
    N528 = 1;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("8. OUTPUT: N545 = %b", N545);
    $display("8. OUTPUT: N1581 = %b", N1581);
    $display("8. OUTPUT: N1901 = %b", N1901);
    $display("8. OUTPUT: N2223 = %b", N2223);
    $display("8. OUTPUT: N2548 = %b", N2548);
    $display("8. OUTPUT: N2877 = %b", N2877);
    $display("8. OUTPUT: N3211 = %b", N3211);
    $display("8. OUTPUT: N3552 = %b", N3552);
    $display("8. OUTPUT: N3895 = %b", N3895);
    $display("8. OUTPUT: N4241 = %b", N4241);
    $display("8. OUTPUT: N4591 = %b", N4591);
    $display("8. OUTPUT: N4946 = %b", N4946);
    $display("8. OUTPUT: N5308 = %b", N5308);
    $display("8. OUTPUT: N5672 = %b", N5672);
    $display("8. OUTPUT: N5971 = %b", N5971);
    $display("8. OUTPUT: N6123 = %b", N6123);
    $display("8. OUTPUT: N6150 = %b", N6150);
    $display("8. OUTPUT: N6160 = %b", N6160);
    $display("8. OUTPUT: N6170 = %b", N6170);
    $display("8. OUTPUT: N6180 = %b", N6180);
    $display("8. OUTPUT: N6190 = %b", N6190);
    $display("8. OUTPUT: N6200 = %b", N6200);
    $display("8. OUTPUT: N6210 = %b", N6210);
    $display("8. OUTPUT: N6220 = %b", N6220);
    $display("8. OUTPUT: N6230 = %b", N6230);
    $display("8. OUTPUT: N6240 = %b", N6240);
    $display("8. OUTPUT: N6250 = %b", N6250);
    $display("8. OUTPUT: N6260 = %b", N6260);
    $display("8. OUTPUT: N6270 = %b", N6270);
    $display("8. OUTPUT: N6280 = %b", N6280);
    $display("8. OUTPUT: N6287 = %b", N6287);
    $display("8. OUTPUT: N6288 = %b", N6288);

    // Aplicando vetor 9
    N1 = 1;
    N18 = 1;
    N35 = 0;
    N52 = 1;
    N69 = 1;
    N86 = 1;
    N103 = 1;
    N120 = 1;
    N137 = 1;
    N154 = 1;
    N171 = 0;
    N188 = 0;
    N205 = 1;
    N222 = 0;
    N239 = 0;
    N256 = 1;
    N273 = 0;
    N290 = 0;
    N307 = 0;
    N324 = 0;
    N341 = 1;
    N358 = 0;
    N375 = 0;
    N392 = 1;
    N409 = 0;
    N426 = 0;
    N443 = 1;
    N460 = 1;
    N477 = 1;
    N494 = 0;
    N511 = 0;
    N528 = 1;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("9. OUTPUT: N545 = %b", N545);
    $display("9. OUTPUT: N1581 = %b", N1581);
    $display("9. OUTPUT: N1901 = %b", N1901);
    $display("9. OUTPUT: N2223 = %b", N2223);
    $display("9. OUTPUT: N2548 = %b", N2548);
    $display("9. OUTPUT: N2877 = %b", N2877);
    $display("9. OUTPUT: N3211 = %b", N3211);
    $display("9. OUTPUT: N3552 = %b", N3552);
    $display("9. OUTPUT: N3895 = %b", N3895);
    $display("9. OUTPUT: N4241 = %b", N4241);
    $display("9. OUTPUT: N4591 = %b", N4591);
    $display("9. OUTPUT: N4946 = %b", N4946);
    $display("9. OUTPUT: N5308 = %b", N5308);
    $display("9. OUTPUT: N5672 = %b", N5672);
    $display("9. OUTPUT: N5971 = %b", N5971);
    $display("9. OUTPUT: N6123 = %b", N6123);
    $display("9. OUTPUT: N6150 = %b", N6150);
    $display("9. OUTPUT: N6160 = %b", N6160);
    $display("9. OUTPUT: N6170 = %b", N6170);
    $display("9. OUTPUT: N6180 = %b", N6180);
    $display("9. OUTPUT: N6190 = %b", N6190);
    $display("9. OUTPUT: N6200 = %b", N6200);
    $display("9. OUTPUT: N6210 = %b", N6210);
    $display("9. OUTPUT: N6220 = %b", N6220);
    $display("9. OUTPUT: N6230 = %b", N6230);
    $display("9. OUTPUT: N6240 = %b", N6240);
    $display("9. OUTPUT: N6250 = %b", N6250);
    $display("9. OUTPUT: N6260 = %b", N6260);
    $display("9. OUTPUT: N6270 = %b", N6270);
    $display("9. OUTPUT: N6280 = %b", N6280);
    $display("9. OUTPUT: N6287 = %b", N6287);
    $display("9. OUTPUT: N6288 = %b", N6288);

    // Aplicando vetor 10
    N1 = 0;
    N18 = 1;
    N35 = 1;
    N52 = 0;
    N69 = 0;
    N86 = 0;
    N103 = 1;
    N120 = 0;
    N137 = 0;
    N154 = 1;
    N171 = 0;
    N188 = 0;
    N205 = 0;
    N222 = 1;
    N239 = 1;
    N256 = 0;
    N273 = 1;
    N290 = 1;
    N307 = 0;
    N324 = 0;
    N341 = 0;
    N358 = 0;
    N375 = 0;
    N392 = 0;
    N409 = 1;
    N426 = 0;
    N443 = 0;
    N460 = 1;
    N477 = 0;
    N494 = 1;
    N511 = 0;
    N528 = 0;

    #5;
    // Falha solicitada sem porta definida; selecionado aleatoriamente 'N2518'
    force uut.N2518 = 1;  // Injetando falha: stuck-at 1 em N2518
    #10;
    $display("10. OUTPUT: N545 = %b", N545);
    $display("10. OUTPUT: N1581 = %b", N1581);
    $display("10. OUTPUT: N1901 = %b", N1901);
    $display("10. OUTPUT: N2223 = %b", N2223);
    $display("10. OUTPUT: N2548 = %b", N2548);
    $display("10. OUTPUT: N2877 = %b", N2877);
    $display("10. OUTPUT: N3211 = %b", N3211);
    $display("10. OUTPUT: N3552 = %b", N3552);
    $display("10. OUTPUT: N3895 = %b", N3895);
    $display("10. OUTPUT: N4241 = %b", N4241);
    $display("10. OUTPUT: N4591 = %b", N4591);
    $display("10. OUTPUT: N4946 = %b", N4946);
    $display("10. OUTPUT: N5308 = %b", N5308);
    $display("10. OUTPUT: N5672 = %b", N5672);
    $display("10. OUTPUT: N5971 = %b", N5971);
    $display("10. OUTPUT: N6123 = %b", N6123);
    $display("10. OUTPUT: N6150 = %b", N6150);
    $display("10. OUTPUT: N6160 = %b", N6160);
    $display("10. OUTPUT: N6170 = %b", N6170);
    $display("10. OUTPUT: N6180 = %b", N6180);
    $display("10. OUTPUT: N6190 = %b", N6190);
    $display("10. OUTPUT: N6200 = %b", N6200);
    $display("10. OUTPUT: N6210 = %b", N6210);
    $display("10. OUTPUT: N6220 = %b", N6220);
    $display("10. OUTPUT: N6230 = %b", N6230);
    $display("10. OUTPUT: N6240 = %b", N6240);
    $display("10. OUTPUT: N6250 = %b", N6250);
    $display("10. OUTPUT: N6260 = %b", N6260);
    $display("10. OUTPUT: N6270 = %b", N6270);
    $display("10. OUTPUT: N6280 = %b", N6280);
    $display("10. OUTPUT: N6287 = %b", N6287);
    $display("10. OUTPUT: N6288 = %b", N6288);

    $finish;
  end
endmodule