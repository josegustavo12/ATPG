module EXEMPLO_AND (input x, input y, output out);
  and u1(out, x, y); // out = x AND y
endmodule